$ full adder example (5.26a)
$ ----------------------------
$(nelist available in page 161 of abramovici text
$ all internal lines are also named in the book)
$
$ 
$ total lines in netlist : 14
$
$
$ 
1gat                   $ ... primary input
2gat                   $ ... primary input
3gat                  $ ... primary input

$
$

11gat		    $ ... primary output
12gat		    $ ... primary output

$
$
$       output         type        inputs
$       ------         ----        ------
        4gat              nand        1gat  2gat
        6gat              nand        1gat  4gat
        7gat              nand        4gat  2gat
        5gat              nand        6gat  7gat
        8gat              nand        3gat 5gat
        9gat              nand        3gat 8gat
        10gat              nand        8gat  5gat
        11gat              nand        9gat  10gat
        12gat             nand        4gat  8gat












		
		
		

